
module WriteBack(clk, rst);
	input wire clk, rst;
endmodule // WriteBack