
module Memory(clk, rst);
	input wire clk, rst;
endmodule // Memory