

module instructionMemory(address, instruction);
	input wire[31:0] address;
	output reg[31:0] instruction;

	always @(*) begin
		case(address/4)
			32'd0: instruction <= 32'b1110_00_1_1101_0_0000_0000_000000010100;
			32'd1: instruction <= 32'b1110_00_1_1101_0_0000_0001_101000000001;
			32'd2: instruction <= 32'b1110_00_1_1101_0_0000_0010_000100000011;
			32'd3: instruction <= 32'b1110_00_0_0100_1_0010_0011_000000000010;
			32'd4: instruction <= 32'b1110_00_0_0101_0_0000_0100_000000000000;
			32'd5: instruction <= 32'b1110_00_0_0010_0_0100_0101_000100000100;
			32'd6: instruction <= 32'b1110_00_0_0110_0_0000_0110_000010100000;
			32'd7: instruction <= 32'b1110_00_0_1100_0_0101_0111_000101000010;
			32'd8: instruction <= 32'b1110_00_0_0000_0_0111_1000_000000000011;
			32'd9: instruction <= 32'b1110_00_0_1111_0_0000_1001_000000000110;
			32'd10: instruction <= 32'b1110_00_0_0001_0_0100_1010_000000000101;
			32'd11: instruction <= 32'b1110_00_0_1010_1_1000_0000_000000000110;
			32'd12: instruction <= 32'b0001_00_0_0100_0_0001_0001_000000000001;
			32'd13: instruction <= 32'b1110_00_0_1000_1_1001_0000_000000001000;
			32'd14: instruction <= 32'b0000_00_0_0100_0_0010_0010_000000000010;
			32'd15: instruction <= 32'b1110_00_1_1101_0_0000_0000_101100000001;
			32'd16: instruction <= 32'b1110_01_0_0100_0_0000_0001_000000000000;
			32'd17: instruction <= 32'b1110_01_0_0100_1_0000_1011_000000000000;
			32'd18: instruction <= 32'b1110_01_0_0100_0_0000_0010_000000000100;
			32'd19: instruction <= 32'b1110_01_0_0100_0_0000_0011_000000001000;
			32'd20: instruction <= 32'b1110_01_0_0100_0_0000_0100_000000001101;
			32'd21: instruction <= 32'b1110_01_0_0100_0_0000_0101_000000010000;
			32'd22: instruction <= 32'b1110_01_0_0100_0_0000_0110_000000010100;
			32'd23: instruction <= 32'b1110_01_0_0100_1_0000_1010_000000000100;
			32'd24: instruction <= 32'b1110_01_0_0100_0_0000_0111_000000011000;
			32'd25: instruction <= 32'b1110_00_1_1101_0_0000_0001_000000000100;
			32'd26: instruction <= 32'b1110_00_1_1101_0_0000_0010_000000000000;
			32'd27: instruction <= 32'b1110_00_1_1101_0_0000_0011_000000000000;
			32'd28: instruction <= 32'b1110_00_0_0100_0_0000_0100_000100000011;
			32'd29: instruction <= 32'b1110_01_0_0100_1_0100_0101_000000000000;
			32'd30: instruction <= 32'b1110_01_0_0100_1_0100_0110_000000000100;
			32'd31: instruction <= 32'b1110_00_0_1010_1_0101_0000_000000000110;
			32'd32: instruction <= 32'b1100_01_0_0100_0_0100_0110_000000000000;
			32'd33: instruction <= 32'b1100_01_0_0100_0_0100_0101_000000000100;
			32'd34: instruction <= 32'b1110_00_1_0100_0_0011_0011_000000000001;
			32'd35: instruction <= 32'b1110_00_1_1010_1_0011_0000_000000000011;
			32'd36: instruction <= 32'b1011_10_1_0_111111111111111111110111;
			32'd37: instruction <= 32'b1110_00_1_0100_0_0010_0010_000000000001;
			32'd38: instruction <= 32'b1110_00_0_1010_1_0010_0000_000000000001;
			32'd39: instruction <= 32'b1011_10_1_0_111111111111111111110010;
			32'd40: instruction <= 32'b1110_01_0_0100_1_0000_0001_000000000000;
			32'd41: instruction <= 32'b1110_01_0_0100_1_0000_0010_000000000100;
			32'd42: instruction <= 32'b1110_01_0_0100_1_0000_0011_000000001000;
			32'd43: instruction <= 32'b1110_01_0_0100_1_0000_0100_000000001100;
			32'd44: instruction <= 32'b1110_01_0_0100_1_0000_0101_000000010000;
			32'd45: instruction <= 32'b1110_01_0_0100_1_0000_0110_000000010100;
			32'd46: instruction <= 32'b1110_10_1_0_111111111111111111111111;
			default: instruction <= 32'd0;
		endcase
	end

endmodule
