
module RegisterUnitMEM2WB(clk, rst);
	input wire clk, rst;
endmodule // RegisterUnitEXE2MEM
