
module RegisterUnitID2EXE(clk, rst);
	input wire clk, rst;
endmodule // RegisterUnitID2EXE
