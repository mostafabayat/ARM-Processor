
module ARM(clk, rst);
	input wire clk, rst;
endmodule // ARM
