
module InstructionDecode(clk, rst);
	input wire clk, rst;
endmodule // ID