
module RegisterUnitEXE2MEM(clk, rst);
	input wire clk, rst;
endmodule // RegisterUnitEXE2MEM
